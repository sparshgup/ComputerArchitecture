`ifndef MEMORY_EXCEPTIONS_H
`define MEMORY_EXCEPTIONS_H

typedef enum logic [2:0] {
  MEM_EXCEPTION_INDEX_MISALIGNED = 0,
  MEM_EXCEPTION_INDEX_OUT_OF_RANGE = 1,
  MEM_EXCEPTION_INDEX_BANK_ERROR = 2,
  MEM_EXCEPTION_INDEX_WRITE_CONFLICT = 3,
  MEM_EXCEPTION_INDEX_READ_WRITE_HAZARD = 4,
  MEM_EXCEPTION_INDEX_MAX
} mem_exception_index_t;

typedef logic [MEM_EXCEPTION_INDEX_MAX-1:0] mem_exception_t;

typedef enum logic [MEM_EXCEPTION_INDEX_MAX-1:0] {
  MEM_EXCEPTION_NONE              = 0,
  MEM_EXCEPTION_MASK_MISALIGNED   = 1 << MEM_EXCEPTION_INDEX_MISALIGNED,
  MEM_EXCEPTION_MASK_OUT_OF_RANGE = 1 << MEM_EXCEPTION_INDEX_OUT_OF_RANGE,
  MEM_EXCEPTION_MASK_BANK_ERROR   = 1 << MEM_EXCEPTION_INDEX_BANK_ERROR,
  MEM_EXCEPTION_MASK_WRITE_CONFLICT = 1 << MEM_EXCEPTION_INDEX_WRITE_CONFLICT,
  MEM_EXCEPTION_MAX_READ_WRITE_HAZARD = 1 << MEM_EXCEPTION_INDEX_READ_WRITE_HAZARD
} mem_exception_mask_t;

`endif // MEMORY_EXCEPTIONS_H
